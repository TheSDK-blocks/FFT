../chisel/verilog/FFT.v